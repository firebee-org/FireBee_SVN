-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 9.1 Build 222 10/21/2009 SJ Full Version"
-- CREATED		"Sat Mar 01 09:20:24 2014"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY firebee1 IS 
	PORT
	(
		FB_ALE :  IN  STD_LOGIC;
		nFB_WR :  IN  STD_LOGIC;
		CLK33M :  IN  STD_LOGIC;
		nFB_CS1 :  IN  STD_LOGIC;
		nFB_CS2 :  IN  STD_LOGIC;
		nFB_CS3 :  IN  STD_LOGIC;
		FB_SIZE0 :  IN  STD_LOGIC;
		FB_SIZE1 :  IN  STD_LOGIC;
		nFB_BURST :  IN  STD_LOGIC;
		LP_BUSY :  IN  STD_LOGIC;
		nACSI_DRQ :  IN  STD_LOGIC;
		nACSI_INT :  IN  STD_LOGIC;
		RxD :  IN  STD_LOGIC;
		CTS :  IN  STD_LOGIC;
		RI :  IN  STD_LOGIC;
		DCD :  IN  STD_LOGIC;
		AMKB_RX :  IN  STD_LOGIC;
		PIC_AMKB_RX :  IN  STD_LOGIC;
		IDE_RDY :  IN  STD_LOGIC;
		IDE_INT :  IN  STD_LOGIC;
		WP_CF_CARD :  IN  STD_LOGIC;
		TRACK00 :  IN  STD_LOGIC;
		nWP :  IN  STD_LOGIC;
		nDCHG :  IN  STD_LOGIC;
		SD_DATA0 :  IN  STD_LOGIC;
		SD_DATA1 :  IN  STD_LOGIC;
		SD_DATA2 :  IN  STD_LOGIC;
		SD_CARD_DEDECT :  IN  STD_LOGIC;
		MIDI_IN :  IN  STD_LOGIC;
		nSCSI_DRQ :  IN  STD_LOGIC;
		SD_WP :  IN  STD_LOGIC;
		nRD_DATA :  IN  STD_LOGIC;
		nSCSI_C_D :  IN  STD_LOGIC;
		nSCSI_I_O :  IN  STD_LOGIC;
		nSCSI_MSG :  IN  STD_LOGIC;
		nDACK0 :  IN  STD_LOGIC;
		PIC_INT :  IN  STD_LOGIC;
		nFB_OE :  IN  STD_LOGIC;
		TOUT0 :  IN  STD_LOGIC;
		nMASTER :  IN  STD_LOGIC;
		DVI_INT :  IN  STD_LOGIC;
		nDACK1 :  IN  STD_LOGIC;
		nPCI_INTD :  IN  STD_LOGIC;
		nPCI_INTC :  IN  STD_LOGIC;
		nPCI_INTB :  IN  STD_LOGIC;
		nPCI_INTA :  IN  STD_LOGIC;
		E0_INT :  IN  STD_LOGIC;
		nINDEX :  IN  STD_LOGIC;
		HD_DD :  IN  STD_LOGIC;
		MAIN_CLK :  IN  STD_LOGIC;
		nRSTO_MCF :  IN  STD_LOGIC;
		SCSI_PAR :  INOUT  STD_LOGIC;
		nSCSI_RST :  INOUT  STD_LOGIC;
		nSCSI_SEL :  INOUT  STD_LOGIC;
		nSCSI_BUSY :  INOUT  STD_LOGIC;
		SD_CD_DATA3 :  INOUT  STD_LOGIC;
		SD_CMD_D1 :  INOUT  STD_LOGIC;
		ACSI_D :  INOUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		FB_AD :  INOUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		IO :  INOUT  STD_LOGIC_VECTOR(17 DOWNTO 0);
		LP_D :  INOUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		SCSI_D :  INOUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		SRD :  INOUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		VD :  INOUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		VDQS :  INOUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		CLK24M576 :  OUT  STD_LOGIC;
		LP_STR :  OUT  STD_LOGIC;
		nACSI_ACK :  OUT  STD_LOGIC;
		nACSI_RESET :  OUT  STD_LOGIC;
		nACSI_CS :  OUT  STD_LOGIC;
		ACSI_DIR :  OUT  STD_LOGIC;
		ACSI_A1 :  OUT  STD_LOGIC;
		nSCSI_ACK :  OUT  STD_LOGIC;
		nSCSI_ATN :  OUT  STD_LOGIC;
		SCSI_DIR :  OUT  STD_LOGIC;
		MIDI_OLR :  OUT  STD_LOGIC;
		MIDI_TLR :  OUT  STD_LOGIC;
		TxD :  OUT  STD_LOGIC;
		RTS :  OUT  STD_LOGIC;
		DTR :  OUT  STD_LOGIC;
		AMKB_TX :  OUT  STD_LOGIC;
		IDE_RES :  OUT  STD_LOGIC;
		nIDE_CS0 :  OUT  STD_LOGIC;
		nIDE_CS1 :  OUT  STD_LOGIC;
		nIDE_WR :  OUT  STD_LOGIC;
		nIDE_RD :  OUT  STD_LOGIC;
		nCF_CS0 :  OUT  STD_LOGIC;
		nCF_CS1 :  OUT  STD_LOGIC;
		nROM3 :  OUT  STD_LOGIC;
		nROM4 :  OUT  STD_LOGIC;
		nRP_UDS :  OUT  STD_LOGIC;
		nRP_LDS :  OUT  STD_LOGIC;
		nSDSEL :  OUT  STD_LOGIC;
		nWR_GATE :  OUT  STD_LOGIC;
		nWR :  OUT  STD_LOGIC;
		YM_QA :  OUT  STD_LOGIC;
		YM_QB :  OUT  STD_LOGIC;
		YM_QC :  OUT  STD_LOGIC;
		SD_CLK :  OUT  STD_LOGIC;
		DSA_D :  OUT  STD_LOGIC;
		nVWE :  OUT  STD_LOGIC;
		nVCAS :  OUT  STD_LOGIC;
		nVRAS :  OUT  STD_LOGIC;
		nVCS :  OUT  STD_LOGIC;
		nPD_VGA :  OUT  STD_LOGIC;
		CLK25M :  OUT  STD_LOGIC;
		TIN0 :  OUT  STD_LOGIC;
		nSRCS :  OUT  STD_LOGIC;
		nSRBLE :  OUT  STD_LOGIC;
		nSRBHE :  OUT  STD_LOGIC;
		nSRWE :  OUT  STD_LOGIC;
		nDREQ1 :  OUT  STD_LOGIC;
		LED_FPGA_OK :  OUT  STD_LOGIC;
		nSROE :  OUT  STD_LOGIC;
		VCKE :  OUT  STD_LOGIC;
		nFB_TA :  OUT  STD_LOGIC;
		nDDR_CLK :  OUT  STD_LOGIC;
		DDR_CLK :  OUT  STD_LOGIC;
		VSYNC_PAD :  OUT  STD_LOGIC;
		HSYNC_PAD :  OUT  STD_LOGIC;
		nBLANK_PAD :  OUT  STD_LOGIC;
		PIXEL_CLK_PAD :  OUT  STD_LOGIC;
		nSYNC :  OUT  STD_LOGIC;
		nMOT_ON :  OUT  STD_LOGIC;
		nSTEP_DIR :  OUT  STD_LOGIC;
		nSTEP :  OUT  STD_LOGIC;
		CLKUSB :  OUT  STD_LOGIC;
		LPDIR :  OUT  STD_LOGIC;
		BA :  OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		nIRQ :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 2);
		VA :  OUT  STD_LOGIC_VECTOR(12 DOWNTO 0);
		VB :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		VDM :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		VG :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		VR :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END firebee1;

ARCHITECTURE bdf_type OF firebee1 IS 

COMPONENT video
	PORT(MAIN_CLK : IN STD_LOGIC;
		 nFB_CS1 : IN STD_LOGIC;
		 nFB_CS2 : IN STD_LOGIC;
		 nFB_CS3 : IN STD_LOGIC;
		 nFB_WR : IN STD_LOGIC;
		 FB_SIZE0 : IN STD_LOGIC;
		 FB_SIZE1 : IN STD_LOGIC;
		 nRSTO : IN STD_LOGIC;
		 nFB_OE : IN STD_LOGIC;
		 FB_ALE : IN STD_LOGIC;
		 DDR_SYNC_66M : IN STD_LOGIC;
		 CLK33M : IN STD_LOGIC;
		 CLK25M : IN STD_LOGIC;
		 CLK_VIDEO : IN STD_LOGIC;
		 VR_BUSY : IN STD_LOGIC;
		 DDRCLK : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 FB_AD : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FB_ADR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 VD : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 VDQS : INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 VR_D : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 VR_RD : OUT STD_LOGIC;
		 nBLANK : OUT STD_LOGIC;
		 nVWE : OUT STD_LOGIC;
		 nVCAS : OUT STD_LOGIC;
		 nVRAS : OUT STD_LOGIC;
		 nVCS : OUT STD_LOGIC;
		 nPD_VGA : OUT STD_LOGIC;
		 VCKE : OUT STD_LOGIC;
		 VSYNC : OUT STD_LOGIC;
		 HSYNC : OUT STD_LOGIC;
		 nSYNC : OUT STD_LOGIC;
		 VIDEO_TA : OUT STD_LOGIC;
		 PIXEL_CLK : OUT STD_LOGIC;
		 VIDEO_RECONFIG : OUT STD_LOGIC;
		 VR_WR : OUT STD_LOGIC;
		 BA : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 VA : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
		 VB : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 VDM : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 VG : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 VR : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT altpll1
	PORT(inclk0 : IN STD_LOGIC;
		 c0 : OUT STD_LOGIC;
		 c1 : OUT STD_LOGIC;
		 c2 : OUT STD_LOGIC;
		 locked : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_ff0
	PORT(clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT altpll2
	PORT(inclk0 : IN STD_LOGIC;
		 c0 : OUT STD_LOGIC;
		 c1 : OUT STD_LOGIC;
		 c2 : OUT STD_LOGIC;
		 c3 : OUT STD_LOGIC;
		 c4 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT altpll3
	PORT(inclk0 : IN STD_LOGIC;
		 c0 : OUT STD_LOGIC;
		 c1 : OUT STD_LOGIC;
		 c2 : OUT STD_LOGIC;
		 c3 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_counter0
	PORT(clock : IN STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
	);
END COMPONENT;

COMPONENT altpll4
	PORT(inclk0 : IN STD_LOGIC;
		 areset : IN STD_LOGIC;
		 scanclk : IN STD_LOGIC;
		 scandata : IN STD_LOGIC;
		 scanclkena : IN STD_LOGIC;
		 configupdate : IN STD_LOGIC;
		 c0 : OUT STD_LOGIC;
		 scandataout : OUT STD_LOGIC;
		 scandone : OUT STD_LOGIC;
		 locked : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT altddio_out3
	PORT(datain_h : IN STD_LOGIC;
		 datain_l : IN STD_LOGIC;
		 outclock : IN STD_LOGIC;
		 dataout : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT altpll_reconfig1
	PORT(reconfig : IN STD_LOGIC;
		 read_param : IN STD_LOGIC;
		 write_param : IN STD_LOGIC;
		 pll_scandataout : IN STD_LOGIC;
		 pll_scandone : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 pll_areset_in : IN STD_LOGIC;
		 counter_param : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 counter_type : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data_in : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 busy : OUT STD_LOGIC;
		 pll_scandata : OUT STD_LOGIC;
		 pll_scanclk : OUT STD_LOGIC;
		 pll_scanclkena : OUT STD_LOGIC;
		 pll_configupdate : OUT STD_LOGIC;
		 pll_areset : OUT STD_LOGIC;
		 data_out : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END COMPONENT;

COMPONENT dsp
	PORT(CLK33M : IN STD_LOGIC;
		 MAIN_CLK : IN STD_LOGIC;
		 nFB_OE : IN STD_LOGIC;
		 nFB_WR : IN STD_LOGIC;
		 nFB_CS1 : IN STD_LOGIC;
		 nFB_CS2 : IN STD_LOGIC;
		 FB_SIZE0 : IN STD_LOGIC;
		 FB_SIZE1 : IN STD_LOGIC;
		 nFB_BURST : IN STD_LOGIC;
		 nRSTO : IN STD_LOGIC;
		 nFB_CS3 : IN STD_LOGIC;
		 FB_AD : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FB_ADR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 IO : INOUT STD_LOGIC_VECTOR(17 DOWNTO 0);
		 SRD : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 nSRCS : OUT STD_LOGIC;
		 nSRBLE : OUT STD_LOGIC;
		 nSRBHE : OUT STD_LOGIC;
		 nSRWE : OUT STD_LOGIC;
		 nSROE : OUT STD_LOGIC;
		 DSP_INT : OUT STD_LOGIC;
		 DSP_TA : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT interrupt_handler
	PORT(MAIN_CLK : IN STD_LOGIC;
		 nFB_WR : IN STD_LOGIC;
		 nFB_CS1 : IN STD_LOGIC;
		 nFB_CS2 : IN STD_LOGIC;
		 FB_SIZE0 : IN STD_LOGIC;
		 FB_SIZE1 : IN STD_LOGIC;
		 PIC_INT : IN STD_LOGIC;
		 E0_INT : IN STD_LOGIC;
		 DVI_INT : IN STD_LOGIC;
		 nPCI_INTA : IN STD_LOGIC;
		 nPCI_INTB : IN STD_LOGIC;
		 nPCI_INTC : IN STD_LOGIC;
		 nPCI_INTD : IN STD_LOGIC;
		 nMFP_INT : IN STD_LOGIC;
		 nFB_OE : IN STD_LOGIC;
		 DSP_INT : IN STD_LOGIC;
		 VSYNC : IN STD_LOGIC;
		 HSYNC : IN STD_LOGIC;
		 DMA_DRQ : IN STD_LOGIC;
		 FB_AD : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FB_ADR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 INT_HANDLER_TA : OUT STD_LOGIC;
		 TIN0 : OUT STD_LOGIC;
		 ACP_CONF : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 nIRQ : OUT STD_LOGIC_VECTOR(7 DOWNTO 2)
	);
END COMPONENT;

COMPONENT falconio_sdcard_ide_cf
	PORT(CLK33M : IN STD_LOGIC;
		 MAIN_CLK : IN STD_LOGIC;
		 CLK2M : IN STD_LOGIC;
		 CLK500k : IN STD_LOGIC;
		 nFB_CS1 : IN STD_LOGIC;
		 FB_SIZE0 : IN STD_LOGIC;
		 FB_SIZE1 : IN STD_LOGIC;
		 nFB_BURST : IN STD_LOGIC;
		 LP_BUSY : IN STD_LOGIC;
		 nACSI_DRQ : IN STD_LOGIC;
		 nACSI_INT : IN STD_LOGIC;
		 nSCSI_DRQ : IN STD_LOGIC;
		 nSCSI_MSG : IN STD_LOGIC;
		 MIDI_IN : IN STD_LOGIC;
		 RxD : IN STD_LOGIC;
		 CTS : IN STD_LOGIC;
		 RI : IN STD_LOGIC;
		 DCD : IN STD_LOGIC;
		 AMKB_RX : IN STD_LOGIC;
		 PIC_AMKB_RX : IN STD_LOGIC;
		 IDE_RDY : IN STD_LOGIC;
		 IDE_INT : IN STD_LOGIC;
		 WP_CS_CARD : IN STD_LOGIC;
		 nINDEX : IN STD_LOGIC;
		 TRACK00 : IN STD_LOGIC;
		 nRD_DATA : IN STD_LOGIC;
		 nDCHG : IN STD_LOGIC;
		 SD_DATA0 : IN STD_LOGIC;
		 SD_DATA1 : IN STD_LOGIC;
		 SD_DATA2 : IN STD_LOGIC;
		 SD_CARD_DEDECT : IN STD_LOGIC;
		 SD_WP : IN STD_LOGIC;
		 nDACK0 : IN STD_LOGIC;
		 nFB_WR : IN STD_LOGIC;
		 WP_CF_CARD : IN STD_LOGIC;
		 nWP : IN STD_LOGIC;
		 nFB_CS2 : IN STD_LOGIC;
		 nRSTO : IN STD_LOGIC;
		 nSCSI_C_D : IN STD_LOGIC;
		 nSCSI_I_O : IN STD_LOGIC;
		 CLK2M4576 : IN STD_LOGIC;
		 nFB_OE : IN STD_LOGIC;
		 VSYNC : IN STD_LOGIC;
		 HSYNC : IN STD_LOGIC;
		 DSP_INT : IN STD_LOGIC;
		 nBLANK : IN STD_LOGIC;
		 FDC_CLK : IN STD_LOGIC;
		 FB_ALE : IN STD_LOGIC;
		 HD_DD : IN STD_LOGIC;
		 SCSI_PAR : INOUT STD_LOGIC;
		 nSCSI_SEL : INOUT STD_LOGIC;
		 nSCSI_BUSY : INOUT STD_LOGIC;
		 nSCSI_RST : INOUT STD_LOGIC;
		 SD_CD_DATA3 : INOUT STD_LOGIC;
		 SD_CDM_D1 : INOUT STD_LOGIC;
		 ACP_CONF : IN STD_LOGIC_VECTOR(31 DOWNTO 24);
		 ACSI_D : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 FB_AD : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FB_ADR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 LP_D : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 SCSI_D : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 nIDE_CS1 : OUT STD_LOGIC;
		 nIDE_CS0 : OUT STD_LOGIC;
		 LP_STR : OUT STD_LOGIC;
		 LP_DIR : OUT STD_LOGIC;
		 nACSI_ACK : OUT STD_LOGIC;
		 nACSI_RESET : OUT STD_LOGIC;
		 nACSI_CS : OUT STD_LOGIC;
		 ACSI_DIR : OUT STD_LOGIC;
		 ACSI_A1 : OUT STD_LOGIC;
		 nSCSI_ACK : OUT STD_LOGIC;
		 nSCSI_ATN : OUT STD_LOGIC;
		 SCSI_DIR : OUT STD_LOGIC;
		 SD_CLK : OUT STD_LOGIC;
		 YM_QA : OUT STD_LOGIC;
		 YM_QC : OUT STD_LOGIC;
		 YM_QB : OUT STD_LOGIC;
		 nSDSEL : OUT STD_LOGIC;
		 STEP : OUT STD_LOGIC;
		 MOT_ON : OUT STD_LOGIC;
		 nRP_LDS : OUT STD_LOGIC;
		 nRP_UDS : OUT STD_LOGIC;
		 nROM4 : OUT STD_LOGIC;
		 nROM3 : OUT STD_LOGIC;
		 nCF_CS1 : OUT STD_LOGIC;
		 nCF_CS0 : OUT STD_LOGIC;
		 nIDE_RD : OUT STD_LOGIC;
		 nIDE_WR : OUT STD_LOGIC;
		 AMKB_TX : OUT STD_LOGIC;
		 IDE_RES : OUT STD_LOGIC;
		 DTR : OUT STD_LOGIC;
		 RTS : OUT STD_LOGIC;
		 TxD : OUT STD_LOGIC;
		 MIDI_OLR : OUT STD_LOGIC;
		 MIDI_TLR : OUT STD_LOGIC;
		 nDREQ0 : OUT STD_LOGIC;
		 DSA_D : OUT STD_LOGIC;
		 nMFP_INT : OUT STD_LOGIC;
		 FALCON_IO_TA : OUT STD_LOGIC;
		 STEP_DIR : OUT STD_LOGIC;
		 WR_DATA : OUT STD_LOGIC;
		 WR_GATE : OUT STD_LOGIC;
		 DMA_DRQ : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	ACP_CONF :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	CLK25M_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	CLK2M :  STD_LOGIC;
SIGNAL	CLK2M4576 :  STD_LOGIC;
SIGNAL	CLK48M :  STD_LOGIC;
SIGNAL	CLK500k :  STD_LOGIC;
SIGNAL	CLK_VIDEO :  STD_LOGIC;
SIGNAL	DDR_SYNC_66M :  STD_LOGIC;
SIGNAL	DDRCLK :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	DMA_DRQ :  STD_LOGIC;
SIGNAL	DSP_INT :  STD_LOGIC;
SIGNAL	DSP_TA :  STD_LOGIC;
SIGNAL	FALCON_IO_TA :  STD_LOGIC;
SIGNAL	FB_ADR :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	FDC_CLK :  STD_LOGIC;
SIGNAL	HSYNC :  STD_LOGIC;
SIGNAL	INT_HANDLER_TA :  STD_LOGIC;
SIGNAL	LP_DIR :  STD_LOGIC;
SIGNAL	MOT_ON :  STD_LOGIC;
SIGNAL	nBLANK :  STD_LOGIC;
SIGNAL	nDREQ0 :  STD_LOGIC;
SIGNAL	nMFP_INT :  STD_LOGIC;
SIGNAL	nRSTO :  STD_LOGIC;
SIGNAL	PIXEL_CLK :  STD_LOGIC;
SIGNAL	SD_CDM_D1 :  STD_LOGIC;
SIGNAL	STEP :  STD_LOGIC;
SIGNAL	STEP_DIR :  STD_LOGIC;
SIGNAL	TIMEBASE :  STD_LOGIC_VECTOR(17 DOWNTO 0);
SIGNAL	VIDEO_RECONFIG :  STD_LOGIC;
SIGNAL	Video_TA :  STD_LOGIC;
SIGNAL	VR_BUSY :  STD_LOGIC;
SIGNAL	VR_D :  STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL	VR_RD :  STD_LOGIC;
SIGNAL	VR_WR :  STD_LOGIC;
SIGNAL	VSYNC :  STD_LOGIC;
SIGNAL	WR_DATA :  STD_LOGIC;
SIGNAL	WR_GATE :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;


BEGIN 
nDREQ1 <= nDACK1;
SYNTHESIZED_WIRE_9 <= '0';
SYNTHESIZED_WIRE_10 <= '1';



b2v_Fredi_Aschwanden : video
PORT MAP(MAIN_CLK => MAIN_CLK,
		 nFB_CS1 => nFB_CS1,
		 nFB_CS2 => nFB_CS2,
		 nFB_CS3 => nFB_CS3,
		 nFB_WR => nFB_WR,
		 FB_SIZE0 => FB_SIZE0,
		 FB_SIZE1 => FB_SIZE1,
		 nRSTO => nRSTO,
		 nFB_OE => nFB_OE,
		 FB_ALE => FB_ALE,
		 DDR_SYNC_66M => DDR_SYNC_66M,
		 CLK33M => CLK33M,
		 CLK25M => CLK25M_ALTERA_SYNTHESIZED,
		 CLK_VIDEO => CLK_VIDEO,
		 VR_BUSY => VR_BUSY,
		 DDRCLK => DDRCLK,
		 FB_AD => FB_AD,
		 FB_ADR => FB_ADR,
		 VD => VD,
		 VDQS => VDQS,
		 VR_D => VR_D,
		 VR_RD => VR_RD,
		 nBLANK => nBLANK,
		 nVWE => nVWE,
		 nVCAS => nVCAS,
		 nVRAS => nVRAS,
		 nVCS => nVCS,
		 nPD_VGA => nPD_VGA,
		 VCKE => VCKE,
		 VSYNC => VSYNC,
		 HSYNC => HSYNC,
		 nSYNC => nSYNC,
		 VIDEO_TA => Video_TA,
		 PIXEL_CLK => PIXEL_CLK,
		 VIDEO_RECONFIG => VIDEO_RECONFIG,
		 VR_WR => VR_WR,
		 BA => BA,
		 VA => VA,
		 VB => VB,
		 VDM => VDM,
		 VG => VG,
		 VR => VR);


b2v_inst : altpll1
PORT MAP(inclk0 => CLK33M,
		 c0 => CLK500k,
		 c1 => CLK2M4576,
		 c2 => CLK24M576,
		 locked => SYNTHESIZED_WIRE_5);


b2v_inst1 : lpm_ff0
PORT MAP(clock => DDR_SYNC_66M,
		 enable => FB_ALE,
		 data => FB_AD,
		 q => FB_ADR);




b2v_inst12 : altpll2
PORT MAP(inclk0 => MAIN_CLK,
		 c0 => DDRCLK(0),
		 c1 => DDRCLK(1),
		 c2 => DDRCLK(2),
		 c3 => DDRCLK(3),
		 c4 => DDR_SYNC_66M);


b2v_inst13 : altpll3
PORT MAP(inclk0 => CLK33M,
		 c0 => CLK2M,
		 c1 => FDC_CLK,
		 c2 => CLK25M_ALTERA_SYNTHESIZED,
		 c3 => CLK48M);


nMOT_ON <= NOT(MOT_ON);



nSTEP_DIR <= NOT(STEP_DIR);



nSTEP <= NOT(STEP);



nWR <= NOT(WR_DATA);



b2v_inst18 : lpm_counter0
PORT MAP(clock => CLK500k,
		 q => TIMEBASE);


nWR_GATE <= NOT(WR_GATE);



nFB_TA <= NOT(Video_TA OR INT_HANDLER_TA OR DSP_TA OR FALCON_IO_TA);


b2v_inst22 : altpll4
PORT MAP(inclk0 => CLK48M,
		 areset => SYNTHESIZED_WIRE_0,
		 scanclk => SYNTHESIZED_WIRE_1,
		 scandata => SYNTHESIZED_WIRE_2,
		 scanclkena => SYNTHESIZED_WIRE_3,
		 configupdate => SYNTHESIZED_WIRE_4,
		 c0 => CLK_VIDEO,
		 scandataout => SYNTHESIZED_WIRE_6,
		 scandone => SYNTHESIZED_WIRE_7);


SYNTHESIZED_WIRE_8 <= NOT(nRSTO);



nRSTO <= SYNTHESIZED_WIRE_5 AND nRSTO_MCF;

LED_FPGA_OK <= TIMEBASE(17);



nDDR_CLK <= NOT(DDRCLK(0));



b2v_inst5 : altddio_out3
PORT MAP(datain_h => VSYNC,
		 datain_l => VSYNC,
		 outclock => PIXEL_CLK,
		 dataout => VSYNC_PAD);


b2v_inst6 : altddio_out3
PORT MAP(datain_h => HSYNC,
		 datain_l => HSYNC,
		 outclock => PIXEL_CLK,
		 dataout => HSYNC_PAD);


b2v_inst7 : altpll_reconfig1
PORT MAP(reconfig => VIDEO_RECONFIG,
		 read_param => VR_RD,
		 write_param => VR_WR,
		 pll_scandataout => SYNTHESIZED_WIRE_6,
		 pll_scandone => SYNTHESIZED_WIRE_7,
		 clock => MAIN_CLK,
		 reset => SYNTHESIZED_WIRE_8,
		 counter_param => FB_ADR(8 DOWNTO 6),
		 counter_type => FB_ADR(5 DOWNTO 2),
		 data_in => FB_AD(24 DOWNTO 16),
		 busy => VR_BUSY,
		 pll_scandata => SYNTHESIZED_WIRE_2,
		 pll_scanclk => SYNTHESIZED_WIRE_1,
		 pll_scanclkena => SYNTHESIZED_WIRE_3,
		 pll_configupdate => SYNTHESIZED_WIRE_4,
		 pll_areset => SYNTHESIZED_WIRE_0,
		 data_out => VR_D);


b2v_inst8 : altddio_out3
PORT MAP(datain_h => nBLANK,
		 datain_l => nBLANK,
		 outclock => PIXEL_CLK,
		 dataout => nBLANK_PAD);


b2v_inst9 : altddio_out3
PORT MAP(datain_h => SYNTHESIZED_WIRE_9,
		 datain_l => SYNTHESIZED_WIRE_10,
		 outclock => PIXEL_CLK,
		 dataout => PIXEL_CLK_PAD);


b2v_Mathias_Alles : dsp
PORT MAP(CLK33M => CLK33M,
		 MAIN_CLK => MAIN_CLK,
		 nFB_OE => nFB_OE,
		 nFB_WR => nFB_WR,
		 nFB_CS1 => nFB_CS1,
		 nFB_CS2 => nFB_CS2,
		 FB_SIZE0 => FB_SIZE0,
		 FB_SIZE1 => FB_SIZE1,
		 nFB_BURST => nFB_BURST,
		 nRSTO => nRSTO,
		 nFB_CS3 => nFB_CS3,
		 FB_AD => FB_AD,
		 FB_ADR => FB_ADR,
		 IO => IO,
		 SRD => SRD,
		 nSRCS => nSRCS,
		 nSRBLE => nSRBLE,
		 nSRBHE => nSRBHE,
		 nSRWE => nSRWE,
		 nSROE => nSROE,
		 DSP_INT => DSP_INT,
		 DSP_TA => DSP_TA);


b2v_nobody : interrupt_handler
PORT MAP(MAIN_CLK => MAIN_CLK,
		 nFB_WR => nFB_WR,
		 nFB_CS1 => nFB_CS1,
		 nFB_CS2 => nFB_CS2,
		 FB_SIZE0 => FB_SIZE0,
		 FB_SIZE1 => FB_SIZE1,
		 PIC_INT => PIC_INT,
		 E0_INT => E0_INT,
		 DVI_INT => DVI_INT,
		 nPCI_INTA => nPCI_INTA,
		 nPCI_INTB => nPCI_INTB,
		 nPCI_INTC => nPCI_INTC,
		 nPCI_INTD => nPCI_INTD,
		 nMFP_INT => nMFP_INT,
		 nFB_OE => nFB_OE,
		 DSP_INT => DSP_INT,
		 VSYNC => VSYNC,
		 HSYNC => HSYNC,
		 DMA_DRQ => DMA_DRQ,
		 FB_AD => FB_AD,
		 FB_ADR => FB_ADR,
		 INT_HANDLER_TA => INT_HANDLER_TA,
		 TIN0 => TIN0,
		 ACP_CONF => ACP_CONF,
		 nIRQ => nIRQ);


b2v_Wolfgang_Foerster_and_Fredi_Aschwanden : falconio_sdcard_ide_cf
PORT MAP(CLK33M => CLK33M,
		 MAIN_CLK => MAIN_CLK,
		 CLK2M => CLK2M,
		 CLK500k => CLK500k,
		 nFB_CS1 => nFB_CS1,
		 FB_SIZE0 => FB_SIZE0,
		 FB_SIZE1 => FB_SIZE1,
		 nFB_BURST => nFB_BURST,
		 LP_BUSY => LP_BUSY,
		 nACSI_DRQ => nACSI_DRQ,
		 nACSI_INT => nACSI_INT,
		 nSCSI_DRQ => nSCSI_DRQ,
		 nSCSI_MSG => nSCSI_MSG,
		 MIDI_IN => MIDI_IN,
		 RxD => RxD,
		 CTS => CTS,
		 RI => RI,
		 DCD => DCD,
		 AMKB_RX => AMKB_RX,
		 PIC_AMKB_RX => PIC_AMKB_RX,
		 IDE_RDY => IDE_RDY,
		 IDE_INT => IDE_INT,
		 nINDEX => nINDEX,
		 TRACK00 => TRACK00,
		 nRD_DATA => nRD_DATA,
		 nDCHG => nDCHG,
		 SD_DATA0 => SD_DATA0,
		 SD_DATA1 => SD_DATA1,
		 SD_DATA2 => SD_DATA2,
		 SD_CARD_DEDECT => SD_CARD_DEDECT,
		 SD_WP => SD_WP,
		 nDACK0 => nDACK0,
		 nFB_WR => nFB_WR,
		 WP_CF_CARD => WP_CF_CARD,
		 nWP => nWP,
		 nFB_CS2 => nFB_CS2,
		 nRSTO => nRSTO,
		 nSCSI_C_D => nSCSI_C_D,
		 nSCSI_I_O => nSCSI_I_O,
		 CLK2M4576 => CLK2M4576,
		 nFB_OE => nFB_OE,
		 VSYNC => VSYNC,
		 HSYNC => HSYNC,
		 DSP_INT => DSP_INT,
		 nBLANK => nBLANK,
		 FDC_CLK => FDC_CLK,
		 FB_ALE => FB_ALE,
		 HD_DD => HD_DD,
		 SCSI_PAR => SCSI_PAR,
		 nSCSI_SEL => nSCSI_SEL,
		 nSCSI_BUSY => nSCSI_BUSY,
		 nSCSI_RST => nSCSI_RST,
		 SD_CD_DATA3 => SD_CD_DATA3,
		 SD_CDM_D1 => SD_CDM_D1,
		 ACP_CONF => ACP_CONF(31 DOWNTO 24),
		 ACSI_D => ACSI_D,
		 FB_AD => FB_AD,
		 FB_ADR => FB_ADR,
		 LP_D => LP_D,
		 SCSI_D => SCSI_D,
		 nIDE_CS1 => nIDE_CS1,
		 nIDE_CS0 => nIDE_CS0,
		 LP_STR => LP_STR,
		 LP_DIR => LP_DIR,
		 nACSI_ACK => nACSI_ACK,
		 nACSI_RESET => nACSI_RESET,
		 nACSI_CS => nACSI_CS,
		 ACSI_DIR => ACSI_DIR,
		 ACSI_A1 => ACSI_A1,
		 nSCSI_ACK => nSCSI_ACK,
		 nSCSI_ATN => nSCSI_ATN,
		 SCSI_DIR => SCSI_DIR,
		 SD_CLK => SD_CLK,
		 YM_QA => YM_QA,
		 YM_QC => YM_QC,
		 YM_QB => YM_QB,
		 nSDSEL => nSDSEL,
		 STEP => STEP,
		 MOT_ON => MOT_ON,
		 nRP_LDS => nRP_LDS,
		 nRP_UDS => nRP_UDS,
		 nROM4 => nROM4,
		 nROM3 => nROM3,
		 nCF_CS1 => nCF_CS1,
		 nCF_CS0 => nCF_CS0,
		 nIDE_RD => nIDE_RD,
		 nIDE_WR => nIDE_WR,
		 AMKB_TX => AMKB_TX,
		 IDE_RES => IDE_RES,
		 DTR => DTR,
		 RTS => RTS,
		 TxD => TxD,
		 MIDI_OLR => MIDI_OLR,
		 MIDI_TLR => MIDI_TLR,
		 DSA_D => DSA_D,
		 nMFP_INT => nMFP_INT,
		 FALCON_IO_TA => FALCON_IO_TA,
		 STEP_DIR => STEP_DIR,
		 WR_DATA => WR_DATA,
		 WR_GATE => WR_GATE,
		 DMA_DRQ => DMA_DRQ);

SD_CMD_D1 <= SD_CDM_D1;
CLK25M <= CLK25M_ALTERA_SYNTHESIZED;
DDR_CLK <= DDRCLK(0);
CLKUSB <= CLK48M;
LPDIR <= LP_DIR;

END bdf_type;