// megafunction wizard: %ALTDDIO_BIDIR%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTDDIO_BIDIR 

// ============================================================
// File Name: altddio_bidir0.v
// Megafunction Name(s):
// 			ALTDDIO_BIDIR
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.1.0 Build 162 10/23/2013 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altddio_bidir0 (
	datain_h,
	datain_l,
	inclock,
	oe,
	outclock,
	combout,
	dataout_h,
	dataout_l,
	padio);

	input	[31:0]  datain_h;
	input	[31:0]  datain_l;
	input	  inclock;
	input	  oe;
	input	  outclock;
	output	[31:0]  combout;
	output	[31:0]  dataout_h;
	output	[31:0]  dataout_l;
	inout	[31:0]  padio;

	wire [31:0] sub_wire0;
	wire [31:0] sub_wire1;
	wire [31:0] sub_wire2;
	wire [31:0] combout = sub_wire0[31:0];
	wire [31:0] dataout_h = sub_wire1[31:0];
	wire [31:0] dataout_l = sub_wire2[31:0];

	altddio_bidir	ALTDDIO_BIDIR_component (
				.padio (padio),
				.datain_h (datain_h),
				.datain_l (datain_l),
				.oe (oe),
				.outclock (outclock),
				.inclock (inclock),
				.combout (sub_wire0),
				.dataout_h (sub_wire1),
				.dataout_l (sub_wire2),
				.aclr (1'b0),
				.aset (1'b0),
				.dqsundelayedout (),
				.inclocken (1'b1),
				.oe_out (),
				.outclocken (1'b1),
				.sclr (1'b0),
				.sset (1'b0));
	defparam
		ALTDDIO_BIDIR_component.extend_oe_disable = "OFF",
		ALTDDIO_BIDIR_component.implement_input_in_lcell = "ON",
		ALTDDIO_BIDIR_component.intended_device_family = "Cyclone III",
		ALTDDIO_BIDIR_component.invert_output = "OFF",
		ALTDDIO_BIDIR_component.lpm_hint = "UNUSED",
		ALTDDIO_BIDIR_component.lpm_type = "altddio_bidir",
		ALTDDIO_BIDIR_component.oe_reg = "UNREGISTERED",
		ALTDDIO_BIDIR_component.power_up_high = "OFF",
		ALTDDIO_BIDIR_component.width = 32;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: CONSTANT: EXTEND_OE_DISABLE STRING "OFF"
// Retrieval info: CONSTANT: IMPLEMENT_INPUT_IN_LCELL STRING "ON"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: CONSTANT: INVERT_OUTPUT STRING "OFF"
// Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altddio_bidir"
// Retrieval info: CONSTANT: OE_REG STRING "UNREGISTERED"
// Retrieval info: CONSTANT: POWER_UP_HIGH STRING "OFF"
// Retrieval info: CONSTANT: WIDTH NUMERIC "32"
// Retrieval info: USED_PORT: combout 0 0 32 0 OUTPUT NODEFVAL "combout[31..0]"
// Retrieval info: CONNECT: combout 0 0 32 0 @combout 0 0 32 0
// Retrieval info: USED_PORT: datain_h 0 0 32 0 INPUT NODEFVAL "datain_h[31..0]"
// Retrieval info: CONNECT: @datain_h 0 0 32 0 datain_h 0 0 32 0
// Retrieval info: USED_PORT: datain_l 0 0 32 0 INPUT NODEFVAL "datain_l[31..0]"
// Retrieval info: CONNECT: @datain_l 0 0 32 0 datain_l 0 0 32 0
// Retrieval info: USED_PORT: dataout_h 0 0 32 0 OUTPUT NODEFVAL "dataout_h[31..0]"
// Retrieval info: CONNECT: dataout_h 0 0 32 0 @dataout_h 0 0 32 0
// Retrieval info: USED_PORT: dataout_l 0 0 32 0 OUTPUT NODEFVAL "dataout_l[31..0]"
// Retrieval info: CONNECT: dataout_l 0 0 32 0 @dataout_l 0 0 32 0
// Retrieval info: USED_PORT: inclock 0 0 0 0 INPUT_CLK_EXT NODEFVAL "inclock"
// Retrieval info: CONNECT: @inclock 0 0 0 0 inclock 0 0 0 0
// Retrieval info: USED_PORT: oe 0 0 0 0 INPUT NODEFVAL "oe"
// Retrieval info: CONNECT: @oe 0 0 0 0 oe 0 0 0 0
// Retrieval info: USED_PORT: outclock 0 0 0 0 INPUT_CLK_EXT NODEFVAL "outclock"
// Retrieval info: CONNECT: @outclock 0 0 0 0 outclock 0 0 0 0
// Retrieval info: USED_PORT: padio 0 0 32 0 BIDIR NODEFVAL "padio[31..0]"
// Retrieval info: CONNECT: padio 0 0 32 0 @padio 0 0 32 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altddio_bidir0.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altddio_bidir0.qip TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altddio_bidir0.bsf FALSE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altddio_bidir0_inst.v FALSE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altddio_bidir0_bb.v FALSE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altddio_bidir0.inc FALSE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altddio_bidir0.cmp FALSE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altddio_bidir0.ppf TRUE FALSE
// Retrieval info: LIB_FILE: altera_mf
