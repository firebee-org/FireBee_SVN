-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 9.1 Build 222 10/21/2009 SJ Full Version"
-- CREATED		"Sat Mar 01 09:19:30 2014"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY video IS 
	PORT
	(
		MAIN_CLK :  IN  STD_LOGIC;
		nFB_CS1 :  IN  STD_LOGIC;
		nFB_CS2 :  IN  STD_LOGIC;
		nFB_CS3 :  IN  STD_LOGIC;
		nFB_WR :  IN  STD_LOGIC;
		FB_SIZE0 :  IN  STD_LOGIC;
		FB_SIZE1 :  IN  STD_LOGIC;
		nRSTO :  IN  STD_LOGIC;
		nFB_OE :  IN  STD_LOGIC;
		FB_ALE :  IN  STD_LOGIC;
		DDR_SYNC_66M :  IN  STD_LOGIC;
		CLK33M :  IN  STD_LOGIC;
		CLK25M :  IN  STD_LOGIC;
		CLK_VIDEO :  IN  STD_LOGIC;
		VR_BUSY :  IN  STD_LOGIC;
		DDRCLK :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		FB_AD :  INOUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		FB_ADR :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		VD :  INOUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		VDQS :  INOUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		VR_D :  IN  STD_LOGIC_VECTOR(8 DOWNTO 0);
		nBLANK :  OUT  STD_LOGIC;
		nVWE :  OUT  STD_LOGIC;
		nVCAS :  OUT  STD_LOGIC;
		nVRAS :  OUT  STD_LOGIC;
		nVCS :  OUT  STD_LOGIC;
		nPD_VGA :  OUT  STD_LOGIC;
		VCKE :  OUT  STD_LOGIC;
		VSYNC :  OUT  STD_LOGIC;
		HSYNC :  OUT  STD_LOGIC;
		nSYNC :  OUT  STD_LOGIC;
		VIDEO_TA :  OUT  STD_LOGIC;
		PIXEL_CLK :  OUT  STD_LOGIC;
		VIDEO_RECONFIG :  OUT  STD_LOGIC;
		VR_WR :  OUT  STD_LOGIC;
		VR_RD :  OUT  STD_LOGIC;
		BA :  OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		VA :  OUT  STD_LOGIC_VECTOR(12 DOWNTO 0);
		VB :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		VDM :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		VG :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		VR :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END video;

ARCHITECTURE bdf_type OF video IS 

ATTRIBUTE black_box : BOOLEAN;
ATTRIBUTE noopt : BOOLEAN;

COMPONENT mux41_0
	PORT(S0 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_0: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_0: COMPONENT IS true;

COMPONENT mux41_1
	PORT(S0 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_1: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_1: COMPONENT IS true;

COMPONENT mux41_2
	PORT(S0 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_2: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_2: COMPONENT IS true;

COMPONENT mux41_3
	PORT(S0 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_3: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_3: COMPONENT IS true;

COMPONENT mux41_4
	PORT(S0 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_4: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_4: COMPONENT IS true;

COMPONENT mux41_5
	PORT(S0 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_5: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_5: COMPONENT IS true;

COMPONENT altdpram2
	PORT(wren_a : IN STD_LOGIC;
		 wren_b : IN STD_LOGIC;
		 clock_a : IN STD_LOGIC;
		 clock_b : IN STD_LOGIC;
		 address_a : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 address_b : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data_a : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data_b : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 q_a : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 q_b : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT blitter
	PORT(nRSTO : IN STD_LOGIC;
		 MAIN_CLK : IN STD_LOGIC;
		 FB_ALE : IN STD_LOGIC;
		 nFB_WR : IN STD_LOGIC;
		 nFB_OE : IN STD_LOGIC;
		 FB_SIZE0 : IN STD_LOGIC;
		 FB_SIZE1 : IN STD_LOGIC;
		 BLITTER_ON : IN STD_LOGIC;
		 nFB_CS1 : IN STD_LOGIC;
		 nFB_CS2 : IN STD_LOGIC;
		 nFB_CS3 : IN STD_LOGIC;
		 DDRCLK0 : IN STD_LOGIC;
		 BLITTER_DACK : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 BLITTER_DIN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 FB_AD : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FB_ADR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 VIDEO_RAM_CTR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 BLITTER_RUN : OUT STD_LOGIC;
		 BLITTER_SIG : OUT STD_LOGIC;
		 BLITTER_WR : OUT STD_LOGIC;
		 BLITTER_TA : OUT STD_LOGIC;
		 BLITTER_ADR : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 BLITTER_DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ddr_ctr
	PORT(nFB_CS1 : IN STD_LOGIC;
		 nFB_CS2 : IN STD_LOGIC;
		 nFB_CS3 : IN STD_LOGIC;
		 nFB_OE : IN STD_LOGIC;
		 FB_SIZE0 : IN STD_LOGIC;
		 FB_SIZE1 : IN STD_LOGIC;
		 nRSTO : IN STD_LOGIC;
		 MAIN_CLK : IN STD_LOGIC;
		 FB_ALE : IN STD_LOGIC;
		 nFB_WR : IN STD_LOGIC;
		 DDR_SYNC_66M : IN STD_LOGIC;
		 BLITTER_SIG : IN STD_LOGIC;
		 BLITTER_WR : IN STD_LOGIC;
		 DDRCLK0 : IN STD_LOGIC;
		 CLK33M : IN STD_LOGIC;
		 CLR_FIFO : IN STD_LOGIC;
		 BLITTER_ADR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FB_AD : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FB_ADR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FIFO_MW : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 VIDEO_RAM_CTR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 nVWE : OUT STD_LOGIC;
		 nVRAS : OUT STD_LOGIC;
		 nVCS : OUT STD_LOGIC;
		 VCKE : OUT STD_LOGIC;
		 nVCAS : OUT STD_LOGIC;
		 SR_FIFO_WRE : OUT STD_LOGIC;
		 SR_DDR_FB : OUT STD_LOGIC;
		 SR_DDR_WR : OUT STD_LOGIC;
		 SR_DDRWR_D_SEL : OUT STD_LOGIC;
		 VIDEO_DDR_TA : OUT STD_LOGIC;
		 SR_BLITTER_DACK : OUT STD_LOGIC;
		 DDRWR_D_SEL1 : OUT STD_LOGIC;
		 BA : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 FB_LE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 FB_VDOE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 SR_VDMP : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 VA : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
		 VDM_SEL : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT altdpram1
	PORT(wren_a : IN STD_LOGIC;
		 wren_b : IN STD_LOGIC;
		 clock_a : IN STD_LOGIC;
		 clock_b : IN STD_LOGIC;
		 address_a : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 address_b : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data_a : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 data_b : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q_a : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q_b : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_fifo_dc0
	PORT(wrreq : IN STD_LOGIC;
		 wrclk : IN STD_LOGIC;
		 rdreq : IN STD_LOGIC;
		 rdclk : IN STD_LOGIC;
		 aclr : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 rdempty : OUT STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		 wrusedw : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END COMPONENT;

COMPONENT altddio_bidir0
	PORT(oe : IN STD_LOGIC;
		 inclock : IN STD_LOGIC;
		 outclock : IN STD_LOGIC;
		 datain_h : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 datain_l : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 padio : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 combout : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 dataout_h : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 dataout_l : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_ff4
	PORT(clock : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_muxvdm
	PORT(data0x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data10x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data11x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data12x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data13x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data14x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data15x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data4x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data5x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data6x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data7x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data8x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data9x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_mux3
	PORT(data1 : IN STD_LOGIC;
		 data0 : IN STD_LOGIC;
		 sel : IN STD_LOGIC;
		 result : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_bustri_long
	PORT(enabledt : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 tridata : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_ff5
	PORT(clock : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_ff1
	PORT(clock : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_ff0
	PORT(clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT altddio_out0
	PORT(outclock : IN STD_LOGIC;
		 datain_h : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 datain_l : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 dataout : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_mux0
	PORT(clock : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_mux5
	PORT(data0x : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_constant2
	PORT(		 result : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_mux1
	PORT(clock : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data4x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data5x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data6x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data7x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_mux2
	PORT(clock : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data10x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data11x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data12x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data13x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data14x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data15x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data4x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data5x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data6x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data7x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data8x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data9x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_shiftreg4
	PORT(clock : IN STD_LOGIC;
		 shiftin : IN STD_LOGIC;
		 shiftout : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_latch0
	PORT(gate : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_ff6
	PORT(clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_ff3
	PORT(clock : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
	);
END COMPONENT;

COMPONENT altddio_out2
	PORT(outclock : IN STD_LOGIC;
		 datain_h : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 datain_l : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 dataout : OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_bustri1
	PORT(enabledt : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 tridata : INOUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_bustri_byt
	PORT(enabledt : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 tridata : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_constant0
	PORT(		 result : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_muxdz
	PORT(clock : IN STD_LOGIC;
		 clken : IN STD_LOGIC;
		 sel : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_fifodz
	PORT(wrreq : IN STD_LOGIC;
		 rdreq : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 aclr : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_bustri3
	PORT(enabledt : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 tridata : INOUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_mux6
	PORT(clock : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 data4x : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 data5x : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 data6x : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 data7x : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_constant1
	PORT(		 result : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_mux4
	PORT(sel : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_constant3
	PORT(		 result : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_shiftreg6
	PORT(clock : IN STD_LOGIC;
		 shiftin : IN STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_shiftreg0
	PORT(load : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 shiftin : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 shiftout : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT altdpram0
	PORT(wren_a : IN STD_LOGIC;
		 wren_b : IN STD_LOGIC;
		 clock_a : IN STD_LOGIC;
		 clock_b : IN STD_LOGIC;
		 address_a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 address_b : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data_a : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 data_b : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 q_a : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 q_b : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END COMPONENT;

COMPONENT video_mod_mux_clutctr
	PORT(nRSTO : IN STD_LOGIC;
		 MAIN_CLK : IN STD_LOGIC;
		 nFB_CS1 : IN STD_LOGIC;
		 nFB_CS2 : IN STD_LOGIC;
		 nFB_CS3 : IN STD_LOGIC;
		 nFB_WR : IN STD_LOGIC;
		 nFB_OE : IN STD_LOGIC;
		 FB_SIZE0 : IN STD_LOGIC;
		 FB_SIZE1 : IN STD_LOGIC;
		 nFB_BURST : IN STD_LOGIC;
		 CLK33M : IN STD_LOGIC;
		 CLK25M : IN STD_LOGIC;
		 BLITTER_RUN : IN STD_LOGIC;
		 CLK_VIDEO : IN STD_LOGIC;
		 VR_BUSY : IN STD_LOGIC;
		 FB_AD : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FB_ADR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 VR_D : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 COLOR8 : OUT STD_LOGIC;
		 ACP_CLUT_RD : OUT STD_LOGIC;
		 COLOR1 : OUT STD_LOGIC;
		 FALCON_CLUT_RDH : OUT STD_LOGIC;
		 FALCON_CLUT_RDL : OUT STD_LOGIC;
		 ST_CLUT_RD : OUT STD_LOGIC;
		 HSYNC : OUT STD_LOGIC;
		 VSYNC : OUT STD_LOGIC;
		 nBLANK : OUT STD_LOGIC;
		 nSYNC : OUT STD_LOGIC;
		 nPD_VGA : OUT STD_LOGIC;
		 FIFO_RDE : OUT STD_LOGIC;
		 COLOR2 : OUT STD_LOGIC;
		 COLOR4 : OUT STD_LOGIC;
		 PIXEL_CLK : OUT STD_LOGIC;
		 BLITTER_ON : OUT STD_LOGIC;
		 VIDEO_MOD_TA : OUT STD_LOGIC;
		 INTER_ZEI : OUT STD_LOGIC;
		 DOP_FIFO_CLR : OUT STD_LOGIC;
		 VIDEO_RECONFIG : OUT STD_LOGIC;
		 VR_WR : OUT STD_LOGIC;
		 VR_RD : OUT STD_LOGIC;
		 CLR_FIFO : OUT STD_LOGIC;
		 ACP_CLUT_WR : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 CCR : OUT STD_LOGIC_VECTOR(23 DOWNTO 0);
		 CCSEL : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 CLUT_MUX_ADR : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 CLUT_OFF : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 FALCON_CLUT_WR : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 ST_CLUT_WR : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 VIDEO_RAM_CTR : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	ACP_CLUT_RD :  STD_LOGIC;
SIGNAL	ACP_CLUT_WR :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	BLITTER_ADR :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BLITTER_DACK :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	BLITTER_DIN :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	BLITTER_DOUT :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	BLITTER_ON :  STD_LOGIC;
SIGNAL	BLITTER_RUN :  STD_LOGIC;
SIGNAL	BLITTER_SIG :  STD_LOGIC;
SIGNAL	BLITTER_TA :  STD_LOGIC;
SIGNAL	BLITTER_WR :  STD_LOGIC;
SIGNAL	CC16 :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	CC24 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	CCA :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	CCF :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	CCR :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	CCS :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	CCSEL :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	CLR_FIFO :  STD_LOGIC;
SIGNAL	CLUT_ADR :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	CLUT_ADR1A :  STD_LOGIC;
SIGNAL	CLUT_ADR2A :  STD_LOGIC;
SIGNAL	CLUT_ADR3A :  STD_LOGIC;
SIGNAL	CLUT_ADR4A :  STD_LOGIC;
SIGNAL	CLUT_ADR5A :  STD_LOGIC;
SIGNAL	CLUT_ADR6A :  STD_LOGIC;
SIGNAL	CLUT_ADR7A :  STD_LOGIC;
SIGNAL	CLUT_MUX_ADR :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	CLUT_OFF :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	COLOR1 :  STD_LOGIC;
SIGNAL	COLOR2 :  STD_LOGIC;
SIGNAL	COLOR4 :  STD_LOGIC;
SIGNAL	COLOR8 :  STD_LOGIC;
SIGNAL	DDR_FB :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	DDR_WR :  STD_LOGIC;
SIGNAL	DDRWR_D_SEL :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	DOP_FIFO_CLR :  STD_LOGIC;
SIGNAL	FALCON_CLUT_RDH :  STD_LOGIC;
SIGNAL	FALCON_CLUT_RDL :  STD_LOGIC;
SIGNAL	FALCON_CLUT_WR :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	FB_DDR :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	FB_LE :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	FB_VDOE :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	FIFO_D :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	FIFO_MW :  STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL	FIFO_RDE :  STD_LOGIC;
SIGNAL	FIFO_WRE :  STD_LOGIC;
SIGNAL	INTER_ZEI :  STD_LOGIC;
SIGNAL	nFB_BURST :  STD_LOGIC;
SIGNAL	PIXEL_CLK_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	SR_BLITTER_DACK :  STD_LOGIC;
SIGNAL	SR_DDR_FB :  STD_LOGIC;
SIGNAL	SR_DDR_WR :  STD_LOGIC;
SIGNAL	SR_DDRWR_D_SEL :  STD_LOGIC;
SIGNAL	SR_FIFO_WRE :  STD_LOGIC;
SIGNAL	SR_VDMP :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	ST_CLUT_RD :  STD_LOGIC;
SIGNAL	ST_CLUT_WR :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	VDM_SEL :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	VDMA :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	VDMB :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	VDMC :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	VDMP :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	VDOUT_OE :  STD_LOGIC;
SIGNAL	VDP_IN :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	VDP_OUT :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	VDR :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	VDVZ :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	VIDEO_DDR_TA :  STD_LOGIC;
SIGNAL	VIDEO_MOD_TA :  STD_LOGIC;
SIGNAL	VIDEO_RAM_CTR :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	ZR_C8 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	ZR_C8B :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	DFF_inst93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	DFF_inst91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC_VECTOR(23 DOWNTO 0);

SIGNAL	GDFX_TEMP_SIGNAL_7 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_8 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_9 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_10 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_11 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_12 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_13 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_14 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_15 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_1 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_2 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_3 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_4 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_5 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_6 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_0 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_16 :  STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN 
VB(7 DOWNTO 0) <= SYNTHESIZED_WIRE_65(7 DOWNTO 0);
VG(7 DOWNTO 0) <= SYNTHESIZED_WIRE_65(15 DOWNTO 8);
VR(7 DOWNTO 0) <= SYNTHESIZED_WIRE_65(23 DOWNTO 16);
SYNTHESIZED_WIRE_0 <= '0';
SYNTHESIZED_WIRE_1 <= '0';
SYNTHESIZED_WIRE_2 <= '0';
SYNTHESIZED_WIRE_3 <= '0';
SYNTHESIZED_WIRE_4 <= '0';
SYNTHESIZED_WIRE_5 <= '0';
SYNTHESIZED_WIRE_19 <= '0';
SYNTHESIZED_WIRE_20 <= '0';
SYNTHESIZED_WIRE_21 <= '0';
SYNTHESIZED_WIRE_22 <= '0';
SYNTHESIZED_WIRE_23 <= '0';
SYNTHESIZED_WIRE_24 <= '0';
SYNTHESIZED_WIRE_55 <= '0';
SYNTHESIZED_WIRE_56 <= '0';
SYNTHESIZED_WIRE_57 <= '0';

GDFX_TEMP_SIGNAL_7 <= (VDMB(119 DOWNTO 0) & VDMA(127 DOWNTO 120));
GDFX_TEMP_SIGNAL_8 <= (VDMB(111 DOWNTO 0) & VDMA(127 DOWNTO 112));
GDFX_TEMP_SIGNAL_9 <= (VDMB(103 DOWNTO 0) & VDMA(127 DOWNTO 104));
GDFX_TEMP_SIGNAL_10 <= (VDMB(95 DOWNTO 0) & VDMA(127 DOWNTO 96));
GDFX_TEMP_SIGNAL_11 <= (VDMB(87 DOWNTO 0) & VDMA(127 DOWNTO 88));
GDFX_TEMP_SIGNAL_12 <= (VDMB(79 DOWNTO 0) & VDMA(127 DOWNTO 80));
GDFX_TEMP_SIGNAL_13 <= (VDMB(71 DOWNTO 0) & VDMA(127 DOWNTO 72));
GDFX_TEMP_SIGNAL_14 <= (VDMB(63 DOWNTO 0) & VDMA(127 DOWNTO 64));
GDFX_TEMP_SIGNAL_15 <= (VDMB(55 DOWNTO 0) & VDMA(127 DOWNTO 56));
GDFX_TEMP_SIGNAL_1 <= (VDMB(47 DOWNTO 0) & VDMA(127 DOWNTO 48));
GDFX_TEMP_SIGNAL_2 <= (VDMB(39 DOWNTO 0) & VDMA(127 DOWNTO 40));
GDFX_TEMP_SIGNAL_3 <= (VDMB(31 DOWNTO 0) & VDMA(127 DOWNTO 32));
GDFX_TEMP_SIGNAL_4 <= (VDMB(23 DOWNTO 0) & VDMA(127 DOWNTO 24));
GDFX_TEMP_SIGNAL_5 <= (VDMB(15 DOWNTO 0) & VDMA(127 DOWNTO 16));
GDFX_TEMP_SIGNAL_6 <= (VDMB(7 DOWNTO 0) & VDMA(127 DOWNTO 8));
CC16(23) <= GDFX_TEMP_SIGNAL_0(15);
CC16(22) <= GDFX_TEMP_SIGNAL_0(14);
CC16(21) <= GDFX_TEMP_SIGNAL_0(13);
CC16(20) <= GDFX_TEMP_SIGNAL_0(12);
CC16(19) <= GDFX_TEMP_SIGNAL_0(11);
CC16(15) <= GDFX_TEMP_SIGNAL_0(10);
CC16(14) <= GDFX_TEMP_SIGNAL_0(9);
CC16(13) <= GDFX_TEMP_SIGNAL_0(8);
CC16(12) <= GDFX_TEMP_SIGNAL_0(7);
CC16(11) <= GDFX_TEMP_SIGNAL_0(6);
CC16(10) <= GDFX_TEMP_SIGNAL_0(5);
CC16(7) <= GDFX_TEMP_SIGNAL_0(4);
CC16(6) <= GDFX_TEMP_SIGNAL_0(3);
CC16(5) <= GDFX_TEMP_SIGNAL_0(2);
CC16(4) <= GDFX_TEMP_SIGNAL_0(1);
CC16(3) <= GDFX_TEMP_SIGNAL_0(0);

CC16(18) <= GDFX_TEMP_SIGNAL_16(7);
CC16(17) <= GDFX_TEMP_SIGNAL_16(6);
CC16(16) <= GDFX_TEMP_SIGNAL_16(5);
CC16(9) <= GDFX_TEMP_SIGNAL_16(4);
CC16(8) <= GDFX_TEMP_SIGNAL_16(3);
CC16(2) <= GDFX_TEMP_SIGNAL_16(2);
CC16(1) <= GDFX_TEMP_SIGNAL_16(1);
CC16(0) <= GDFX_TEMP_SIGNAL_16(0);



b2v_ACP_CLUT_RAM : altdpram2
PORT MAP(wren_a => ACP_CLUT_WR(3),
		 wren_b => SYNTHESIZED_WIRE_0,
		 clock_a => MAIN_CLK,
		 clock_b => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 address_a => FB_ADR(9 DOWNTO 2),
		 address_b => ZR_C8B,
		 data_a => FB_AD(7 DOWNTO 0),
		 q_a => SYNTHESIZED_WIRE_30,
		 q_b => CCA(7 DOWNTO 0));


b2v_ACP_CLUT_RAM54 : altdpram2
PORT MAP(wren_a => ACP_CLUT_WR(2),
		 wren_b => SYNTHESIZED_WIRE_1,
		 clock_a => MAIN_CLK,
		 clock_b => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 address_a => FB_ADR(9 DOWNTO 2),
		 address_b => ZR_C8B,
		 data_a => FB_AD(15 DOWNTO 8),
		 q_a => SYNTHESIZED_WIRE_32,
		 q_b => CCA(15 DOWNTO 8));


b2v_ACP_CLUT_RAM55 : altdpram2
PORT MAP(wren_a => ACP_CLUT_WR(1),
		 wren_b => SYNTHESIZED_WIRE_2,
		 clock_a => MAIN_CLK,
		 clock_b => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 address_a => FB_ADR(9 DOWNTO 2),
		 address_b => ZR_C8B,
		 data_a => FB_AD(23 DOWNTO 16),
		 q_a => SYNTHESIZED_WIRE_33,
		 q_b => CCA(23 DOWNTO 16));


b2v_BLITTER : blitter
PORT MAP(nRSTO => nRSTO,
		 MAIN_CLK => MAIN_CLK,
		 FB_ALE => FB_ALE,
		 nFB_WR => nFB_WR,
		 nFB_OE => nFB_OE,
		 FB_SIZE0 => FB_SIZE0,
		 FB_SIZE1 => FB_SIZE1,
		 BLITTER_ON => BLITTER_ON,
		 nFB_CS1 => nFB_CS1,
		 nFB_CS2 => nFB_CS2,
		 nFB_CS3 => nFB_CS3,
		 DDRCLK0 => DDRCLK(0),
		 BLITTER_DACK => BLITTER_DACK,
		 BLITTER_DIN => BLITTER_DIN,
		 FB_AD => FB_AD,
		 FB_ADR => FB_ADR,
		 VIDEO_RAM_CTR => VIDEO_RAM_CTR,
		 BLITTER_RUN => BLITTER_RUN,
		 BLITTER_SIG => BLITTER_SIG,
		 BLITTER_WR => BLITTER_WR,
		 BLITTER_TA => BLITTER_TA,
		 BLITTER_ADR => BLITTER_ADR,
		 BLITTER_DOUT => BLITTER_DOUT);


b2v_DDR_CTR : ddr_ctr
PORT MAP(nFB_CS1 => nFB_CS1,
		 nFB_CS2 => nFB_CS2,
		 nFB_CS3 => nFB_CS3,
		 nFB_OE => nFB_OE,
		 FB_SIZE0 => FB_SIZE0,
		 FB_SIZE1 => FB_SIZE1,
		 nRSTO => nRSTO,
		 MAIN_CLK => MAIN_CLK,
		 FB_ALE => FB_ALE,
		 nFB_WR => nFB_WR,
		 DDR_SYNC_66M => DDR_SYNC_66M,
		 BLITTER_SIG => BLITTER_SIG,
		 BLITTER_WR => BLITTER_WR,
		 DDRCLK0 => DDRCLK(0),
		 CLK33M => CLK33M,
		 CLR_FIFO => CLR_FIFO,
		 BLITTER_ADR => BLITTER_ADR,
		 FB_AD => FB_AD,
		 FB_ADR => FB_ADR,
		 FIFO_MW => FIFO_MW,
		 VIDEO_RAM_CTR => VIDEO_RAM_CTR,
		 nVWE => nVWE,
		 nVRAS => nVRAS,
		 nVCS => nVCS,
		 VCKE => VCKE,
		 nVCAS => nVCAS,
		 SR_FIFO_WRE => SR_FIFO_WRE,
		 SR_DDR_FB => SR_DDR_FB,
		 SR_DDR_WR => SR_DDR_WR,
		 SR_DDRWR_D_SEL => SR_DDRWR_D_SEL,
		 VIDEO_DDR_TA => VIDEO_DDR_TA,
		 SR_BLITTER_DACK => SR_BLITTER_DACK,
		 DDRWR_D_SEL1 => DDRWR_D_SEL(1),
		 BA => BA,
		 FB_LE => FB_LE,
		 FB_VDOE => FB_VDOE,
		 SR_VDMP => SR_VDMP,
		 VA => VA,
		 VDM_SEL => VDM_SEL);


b2v_FALCON_CLUT_BLUE : altdpram1
PORT MAP(wren_a => FALCON_CLUT_WR(3),
		 wren_b => SYNTHESIZED_WIRE_3,
		 clock_a => MAIN_CLK,
		 clock_b => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 address_a => FB_ADR(9 DOWNTO 2),
		 address_b => CLUT_ADR,
		 data_a => FB_AD(23 DOWNTO 18),
		 q_a => SYNTHESIZED_WIRE_45,
		 q_b => CCF(7 DOWNTO 2));


b2v_FALCON_CLUT_GREEN : altdpram1
PORT MAP(wren_a => FALCON_CLUT_WR(1),
		 wren_b => SYNTHESIZED_WIRE_4,
		 clock_a => MAIN_CLK,
		 clock_b => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 address_a => FB_ADR(9 DOWNTO 2),
		 address_b => CLUT_ADR,
		 data_a => FB_AD(23 DOWNTO 18),
		 q_a => SYNTHESIZED_WIRE_44,
		 q_b => CCF(15 DOWNTO 10));


b2v_FALCON_CLUT_RED : altdpram1
PORT MAP(wren_a => FALCON_CLUT_WR(0),
		 wren_b => SYNTHESIZED_WIRE_5,
		 clock_a => MAIN_CLK,
		 clock_b => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 address_a => FB_ADR(9 DOWNTO 2),
		 address_b => CLUT_ADR,
		 data_a => FB_AD(31 DOWNTO 26),
		 q_a => SYNTHESIZED_WIRE_41,
		 q_b => CCF(23 DOWNTO 18));


b2v_inst : lpm_fifo_dc0
PORT MAP(wrreq => FIFO_WRE,
		 wrclk => DDRCLK(0),
		 rdreq => SYNTHESIZED_WIRE_60,
		 rdclk => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 aclr => CLR_FIFO,
		 data => VDMC,
		 q => SYNTHESIZED_WIRE_63,
		 wrusedw => FIFO_MW);


b2v_inst1 : altddio_bidir0
PORT MAP(oe => VDOUT_OE,
		 inclock => DDRCLK(1),
		 outclock => DDRCLK(3),
		 datain_h => VDP_OUT(63 DOWNTO 32),
		 datain_l => VDP_OUT(31 DOWNTO 0),
		 padio => VD,
		 combout => SYNTHESIZED_WIRE_15,
		 dataout_h => VDP_IN(31 DOWNTO 0),
		 dataout_l => VDP_IN(63 DOWNTO 32));


b2v_inst10 : lpm_ff4
PORT MAP(clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 data => SYNTHESIZED_WIRE_7,
		 q => GDFX_TEMP_SIGNAL_0);


b2v_inst100 : lpm_muxvdm
PORT MAP(data0x => VDMB,
		 data10x => GDFX_TEMP_SIGNAL_1,
		 data11x => GDFX_TEMP_SIGNAL_2,
		 data12x => GDFX_TEMP_SIGNAL_3,
		 data13x => GDFX_TEMP_SIGNAL_4,
		 data14x => GDFX_TEMP_SIGNAL_5,
		 data15x => GDFX_TEMP_SIGNAL_6,
		 data1x => GDFX_TEMP_SIGNAL_7,
		 data2x => GDFX_TEMP_SIGNAL_8,
		 data3x => GDFX_TEMP_SIGNAL_9,
		 data4x => GDFX_TEMP_SIGNAL_10,
		 data5x => GDFX_TEMP_SIGNAL_11,
		 data6x => GDFX_TEMP_SIGNAL_12,
		 data7x => GDFX_TEMP_SIGNAL_13,
		 data8x => GDFX_TEMP_SIGNAL_14,
		 data9x => GDFX_TEMP_SIGNAL_15,
		 sel => VDM_SEL,
		 result => VDMC);


b2v_inst102 : lpm_mux3
PORT MAP(data1 => DFF_inst93,
		 data0 => ZR_C8(0),
		 sel => COLOR1,
		 result => ZR_C8B(0));


CLUT_ADR(4) <= CLUT_OFF(0) OR SYNTHESIZED_WIRE_8;


CLUT_ADR(6) <= CLUT_OFF(2) OR SYNTHESIZED_WIRE_9;


SYNTHESIZED_WIRE_61 <= COLOR8 OR COLOR4;


CLUT_ADR(2) <= CLUT_ADR2A AND SYNTHESIZED_WIRE_61;


SYNTHESIZED_WIRE_16 <= COLOR4 OR COLOR8 OR COLOR2;


b2v_inst108 : lpm_bustri_long
PORT MAP(enabledt => FB_VDOE(0),
		 data => VDR,
		 tridata => FB_AD);


b2v_inst109 : lpm_bustri_long
PORT MAP(enabledt => FB_VDOE(1),
		 data => SYNTHESIZED_WIRE_11,
		 tridata => FB_AD);


b2v_inst11 : lpm_ff5
PORT MAP(clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 data => SYNTHESIZED_WIRE_12,
		 q => ZR_C8);


b2v_inst110 : lpm_bustri_long
PORT MAP(enabledt => FB_VDOE(2),
		 data => SYNTHESIZED_WIRE_13,
		 tridata => FB_AD);


b2v_inst119 : lpm_bustri_long
PORT MAP(enabledt => FB_VDOE(3),
		 data => SYNTHESIZED_WIRE_14,
		 tridata => FB_AD);


b2v_inst12 : lpm_ff1
PORT MAP(clock => DDRCLK(0),
		 data => VDP_IN(31 DOWNTO 0),
		 q => VDVZ(31 DOWNTO 0));


b2v_inst13 : lpm_ff0
PORT MAP(clock => DDR_SYNC_66M,
		 enable => FB_LE(0),
		 data => FB_AD,
		 q => FB_DDR(127 DOWNTO 96));


b2v_inst14 : lpm_ff0
PORT MAP(clock => DDR_SYNC_66M,
		 enable => FB_LE(1),
		 data => FB_AD,
		 q => FB_DDR(95 DOWNTO 64));


b2v_inst15 : lpm_ff0
PORT MAP(clock => DDR_SYNC_66M,
		 enable => FB_LE(2),
		 data => FB_AD,
		 q => FB_DDR(63 DOWNTO 32));


b2v_inst16 : lpm_ff0
PORT MAP(clock => DDR_SYNC_66M,
		 enable => FB_LE(3),
		 data => FB_AD,
		 q => FB_DDR(31 DOWNTO 0));


b2v_inst17 : lpm_ff0
PORT MAP(clock => DDRCLK(0),
		 enable => DDR_FB(1),
		 data => VDP_IN(31 DOWNTO 0),
		 q => SYNTHESIZED_WIRE_11);


b2v_inst18 : lpm_ff0
PORT MAP(clock => DDRCLK(0),
		 enable => DDR_FB(0),
		 data => VDP_IN(63 DOWNTO 32),
		 q => SYNTHESIZED_WIRE_13);


b2v_inst19 : lpm_ff0
PORT MAP(clock => DDRCLK(0),
		 enable => DDR_FB(0),
		 data => VDP_IN(31 DOWNTO 0),
		 q => SYNTHESIZED_WIRE_14);


b2v_inst2 : altddio_out0
PORT MAP(outclock => DDRCLK(3),
		 datain_h => VDMP(7 DOWNTO 4),
		 datain_l => VDMP(3 DOWNTO 0),
		 dataout => VDM);


b2v_inst20 : lpm_ff1
PORT MAP(clock => DDRCLK(0),
		 data => VDVZ(31 DOWNTO 0),
		 q => VDVZ(95 DOWNTO 64));


b2v_inst21 : lpm_mux0
PORT MAP(clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 data0x => FIFO_D(127 DOWNTO 96),
		 data1x => FIFO_D(95 DOWNTO 64),
		 data2x => FIFO_D(63 DOWNTO 32),
		 data3x => FIFO_D(31 DOWNTO 0),
		 sel => CLUT_MUX_ADR(1 DOWNTO 0),
		 result => SYNTHESIZED_WIRE_48);


b2v_inst22 : lpm_mux5
PORT MAP(data0x => FB_DDR(127 DOWNTO 64),
		 data1x => FB_DDR(63 DOWNTO 0),
		 data2x => BLITTER_DOUT(127 DOWNTO 64),
		 data3x => BLITTER_DOUT(63 DOWNTO 0),
		 sel => DDRWR_D_SEL,
		 result => VDP_OUT);


b2v_inst23 : lpm_constant2
PORT MAP(		 result => GDFX_TEMP_SIGNAL_16);


b2v_inst24 : lpm_mux1
PORT MAP(clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 data0x => FIFO_D(127 DOWNTO 112),
		 data1x => FIFO_D(111 DOWNTO 96),
		 data2x => FIFO_D(95 DOWNTO 80),
		 data3x => FIFO_D(79 DOWNTO 64),
		 data4x => FIFO_D(63 DOWNTO 48),
		 data5x => FIFO_D(47 DOWNTO 32),
		 data6x => FIFO_D(31 DOWNTO 16),
		 data7x => FIFO_D(15 DOWNTO 0),
		 sel => CLUT_MUX_ADR(2 DOWNTO 0),
		 result => SYNTHESIZED_WIRE_7);


b2v_inst25 : lpm_mux2
PORT MAP(clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 data0x => FIFO_D(127 DOWNTO 120),
		 data10x => FIFO_D(47 DOWNTO 40),
		 data11x => FIFO_D(39 DOWNTO 32),
		 data12x => FIFO_D(31 DOWNTO 24),
		 data13x => FIFO_D(23 DOWNTO 16),
		 data14x => FIFO_D(15 DOWNTO 8),
		 data15x => FIFO_D(7 DOWNTO 0),
		 data1x => FIFO_D(119 DOWNTO 112),
		 data2x => FIFO_D(111 DOWNTO 104),
		 data3x => FIFO_D(103 DOWNTO 96),
		 data4x => FIFO_D(95 DOWNTO 88),
		 data5x => FIFO_D(87 DOWNTO 80),
		 data6x => FIFO_D(79 DOWNTO 72),
		 data7x => FIFO_D(71 DOWNTO 64),
		 data8x => FIFO_D(63 DOWNTO 56),
		 data9x => FIFO_D(55 DOWNTO 48),
		 sel => CLUT_MUX_ADR,
		 result => SYNTHESIZED_WIRE_12);


b2v_inst26 : lpm_shiftreg4
PORT MAP(clock => DDRCLK(0),
		 shiftin => SR_FIFO_WRE,
		 shiftout => FIFO_WRE);


b2v_inst27 : lpm_latch0
PORT MAP(gate => DDR_SYNC_66M,
		 data => SYNTHESIZED_WIRE_15,
		 q => VDR);



CLUT_ADR(1) <= CLUT_ADR1A AND SYNTHESIZED_WIRE_16;


b2v_inst3 : lpm_ff1
PORT MAP(clock => DDRCLK(0),
		 data => VDP_IN(63 DOWNTO 32),
		 q => VDVZ(63 DOWNTO 32));


CLUT_ADR(3) <= SYNTHESIZED_WIRE_61 AND CLUT_ADR3A;


CLUT_ADR(5) <= CLUT_OFF(1) OR SYNTHESIZED_WIRE_18;


SYNTHESIZED_WIRE_8 <= CLUT_ADR4A AND COLOR8;


SYNTHESIZED_WIRE_18 <= CLUT_ADR5A AND COLOR8;


SYNTHESIZED_WIRE_9 <= CLUT_ADR6A AND COLOR8;


SYNTHESIZED_WIRE_46 <= CLUT_ADR7A AND COLOR8;


b2v_inst36 : lpm_ff6
PORT MAP(clock => DDRCLK(0),
		 enable => BLITTER_DACK(0),
		 data => VDVZ,
		 q => BLITTER_DIN);


VDOUT_OE <= DDR_WR OR SR_DDR_WR;



VIDEO_TA <= BLITTER_TA OR VIDEO_MOD_TA OR VIDEO_DDR_TA;


b2v_inst4 : lpm_ff1
PORT MAP(clock => DDRCLK(0),
		 data => VDVZ(63 DOWNTO 32),
		 q => VDVZ(127 DOWNTO 96));


b2v_inst40 : mux41_0
PORT MAP(S0 => COLOR2,
		 S1 => COLOR4,
		 D0 => CLUT_ADR6A,
		 INH => SYNTHESIZED_WIRE_19,
		 D1 => CLUT_ADR7A,
		 Q => SYNTHESIZED_WIRE_54);


b2v_inst41 : mux41_1
PORT MAP(S0 => COLOR2,
		 S1 => COLOR4,
		 D0 => CLUT_ADR5A,
		 INH => SYNTHESIZED_WIRE_20,
		 D1 => CLUT_ADR6A,
		 Q => SYNTHESIZED_WIRE_53);


b2v_inst42 : mux41_2
PORT MAP(S0 => COLOR2,
		 D2 => CLUT_ADR7A,
		 S1 => COLOR4,
		 D0 => CLUT_ADR4A,
		 INH => SYNTHESIZED_WIRE_21,
		 D1 => CLUT_ADR5A,
		 Q => SYNTHESIZED_WIRE_52);


b2v_inst43 : mux41_3
PORT MAP(S0 => COLOR2,
		 D2 => CLUT_ADR6A,
		 S1 => COLOR4,
		 D0 => CLUT_ADR3A,
		 INH => SYNTHESIZED_WIRE_22,
		 D1 => CLUT_ADR4A,
		 Q => SYNTHESIZED_WIRE_51);


b2v_inst44 : mux41_4
PORT MAP(S0 => COLOR2,
		 D2 => CLUT_ADR5A,
		 S1 => COLOR4,
		 D0 => CLUT_ADR2A,
		 INH => SYNTHESIZED_WIRE_23,
		 D1 => CLUT_ADR3A,
		 Q => SYNTHESIZED_WIRE_50);


b2v_inst45 : mux41_5
PORT MAP(S0 => COLOR2,
		 D2 => CLUT_ADR4A,
		 S1 => COLOR4,
		 D0 => CLUT_ADR1A,
		 INH => SYNTHESIZED_WIRE_24,
		 D1 => CLUT_ADR2A,
		 Q => SYNTHESIZED_WIRE_49);


b2v_inst46 : lpm_ff3
PORT MAP(clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 data => SYNTHESIZED_WIRE_25,
		 q => SYNTHESIZED_WIRE_43);


b2v_inst47 : lpm_ff3
PORT MAP(clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 data => CCF,
		 q => SYNTHESIZED_WIRE_25);



b2v_inst49 : lpm_ff3
PORT MAP(clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 data => SYNTHESIZED_WIRE_26,
		 q => SYNTHESIZED_WIRE_42);


b2v_inst5 : altddio_out2
PORT MAP(outclock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 datain_h => SYNTHESIZED_WIRE_62,
		 datain_l => SYNTHESIZED_WIRE_62,
		 dataout => SYNTHESIZED_WIRE_65);



b2v_inst51 : lpm_bustri1
PORT MAP(enabledt => ST_CLUT_RD,
		 data => SYNTHESIZED_WIRE_29,
		 tridata => FB_AD(26 DOWNTO 24));


b2v_inst52 : lpm_ff3
PORT MAP(clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 data => CCS,
		 q => SYNTHESIZED_WIRE_26);


b2v_inst53 : lpm_bustri_byt
PORT MAP(enabledt => ACP_CLUT_RD,
		 data => SYNTHESIZED_WIRE_30,
		 tridata => FB_AD(7 DOWNTO 0));


b2v_inst54 : lpm_constant0
PORT MAP(		 result => CCS(20 DOWNTO 16));



b2v_inst56 : lpm_bustri1
PORT MAP(enabledt => ST_CLUT_RD,
		 data => SYNTHESIZED_WIRE_31,
		 tridata => FB_AD(22 DOWNTO 20));


b2v_inst57 : lpm_bustri_byt
PORT MAP(enabledt => ACP_CLUT_RD,
		 data => SYNTHESIZED_WIRE_32,
		 tridata => FB_AD(15 DOWNTO 8));


b2v_inst58 : lpm_bustri_byt
PORT MAP(enabledt => ACP_CLUT_RD,
		 data => SYNTHESIZED_WIRE_33,
		 tridata => FB_AD(23 DOWNTO 16));


b2v_inst59 : lpm_constant0
PORT MAP(		 result => CCS(12 DOWNTO 8));




b2v_inst61 : lpm_bustri1
PORT MAP(enabledt => ST_CLUT_RD,
		 data => SYNTHESIZED_WIRE_34,
		 tridata => FB_AD(18 DOWNTO 16));


b2v_inst62 : lpm_muxdz
PORT MAP(clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 clken => FIFO_RDE,
		 sel => INTER_ZEI,
		 data0x => SYNTHESIZED_WIRE_63,
		 data1x => SYNTHESIZED_WIRE_36,
		 result => FIFO_D);


b2v_inst63 : lpm_fifodz
PORT MAP(wrreq => SYNTHESIZED_WIRE_60,
		 rdreq => SYNTHESIZED_WIRE_38,
		 clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 aclr => DOP_FIFO_CLR,
		 data => SYNTHESIZED_WIRE_63,
		 q => SYNTHESIZED_WIRE_36);


b2v_inst64 : lpm_constant0
PORT MAP(		 result => CCS(4 DOWNTO 0));


SYNTHESIZED_WIRE_60 <= FIFO_RDE AND SYNTHESIZED_WIRE_40;


b2v_inst66 : lpm_bustri3
PORT MAP(enabledt => FALCON_CLUT_RDH,
		 data => SYNTHESIZED_WIRE_41,
		 tridata => FB_AD(31 DOWNTO 26));


SYNTHESIZED_WIRE_38 <= FIFO_RDE AND INTER_ZEI;



SYNTHESIZED_WIRE_40 <= NOT(INTER_ZEI);



b2v_inst7 : lpm_mux6
PORT MAP(clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 data0x => SYNTHESIZED_WIRE_42,
		 data1x => SYNTHESIZED_WIRE_43,
		 data4x => CCA,
		 data5x => CC16,
		 data6x => CC24(23 DOWNTO 0),
		 data7x => CCR,
		 sel => CCSEL,
		 result => SYNTHESIZED_WIRE_62);


b2v_inst70 : lpm_bustri3
PORT MAP(enabledt => FALCON_CLUT_RDH,
		 data => SYNTHESIZED_WIRE_44,
		 tridata => FB_AD(23 DOWNTO 18));


b2v_inst71 : lpm_ff6
PORT MAP(clock => DDRCLK(0),
		 enable => FIFO_WRE,
		 data => VDVZ,
		 q => VDMA);




b2v_inst74 : lpm_bustri3
PORT MAP(enabledt => FALCON_CLUT_RDL,
		 data => SYNTHESIZED_WIRE_45,
		 tridata => FB_AD(23 DOWNTO 18));




b2v_inst77 : lpm_constant1
PORT MAP(		 result => CCF(1 DOWNTO 0));



CLUT_ADR(7) <= CLUT_OFF(3) OR SYNTHESIZED_WIRE_46;



b2v_inst80 : lpm_constant1
PORT MAP(		 result => CCF(9 DOWNTO 8));


b2v_inst81 : lpm_mux4
PORT MAP(sel => COLOR1,
		 data0x => ZR_C8(7 DOWNTO 1),
		 data1x => SYNTHESIZED_WIRE_47,
		 result => ZR_C8B(7 DOWNTO 1));


b2v_inst82 : lpm_constant3
PORT MAP(		 result => SYNTHESIZED_WIRE_47);


b2v_inst83 : lpm_constant1
PORT MAP(		 result => CCF(17 DOWNTO 16));


PROCESS(DDRCLK(0),DDR_WR)
BEGIN
if (DDR_WR = '1') THEN
	VDQS(3) <= DDRCLK(0);
ELSE
	VDQS(3) <= 'Z';
END IF;
END PROCESS;


PROCESS(DDRCLK(0),DDR_WR)
BEGIN
if (DDR_WR = '1') THEN
	VDQS(2) <= DDRCLK(0);
ELSE
	VDQS(2) <= 'Z';
END IF;
END PROCESS;


PROCESS(DDRCLK(0),DDR_WR)
BEGIN
if (DDR_WR = '1') THEN
	VDQS(1) <= DDRCLK(0);
ELSE
	VDQS(1) <= 'Z';
END IF;
END PROCESS;


PROCESS(DDRCLK(0),DDR_WR)
BEGIN
if (DDR_WR = '1') THEN
	VDQS(0) <= DDRCLK(0);
ELSE
	VDQS(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(DDRCLK(3))
BEGIN
IF (RISING_EDGE(DDRCLK(3))) THEN
	DDRWR_D_SEL(0) <= SR_DDRWR_D_SEL;
END IF;
END PROCESS;


b2v_inst89 : lpm_shiftreg6
PORT MAP(clock => DDRCLK(0),
		 shiftin => SR_BLITTER_DACK,
		 q => BLITTER_DACK);


b2v_inst9 : lpm_ff1
PORT MAP(clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 data => SYNTHESIZED_WIRE_48,
		 q => CC24);


PROCESS(DDRCLK(3))
BEGIN
IF (RISING_EDGE(DDRCLK(3))) THEN
	DDR_WR <= SR_DDR_WR;
END IF;
END PROCESS;


PROCESS(PIXEL_CLK_ALTERA_SYNTHESIZED)
BEGIN
IF (RISING_EDGE(PIXEL_CLK_ALTERA_SYNTHESIZED)) THEN
	DFF_inst91 <= CLUT_ADR(0);
END IF;
END PROCESS;


b2v_inst92 : lpm_shiftreg6
PORT MAP(clock => DDRCLK(0),
		 shiftin => SR_DDR_FB,
		 q => DDR_FB);


PROCESS(PIXEL_CLK_ALTERA_SYNTHESIZED)
BEGIN
IF (RISING_EDGE(PIXEL_CLK_ALTERA_SYNTHESIZED)) THEN
	DFF_inst93 <= DFF_inst91;
END IF;
END PROCESS;


b2v_inst94 : lpm_ff6
PORT MAP(clock => DDRCLK(0),
		 enable => FIFO_WRE,
		 data => VDMA,
		 q => VDMB);


PROCESS(PIXEL_CLK_ALTERA_SYNTHESIZED)
BEGIN
IF (RISING_EDGE(PIXEL_CLK_ALTERA_SYNTHESIZED)) THEN
	SYNTHESIZED_WIRE_64 <= FIFO_RDE;
END IF;
END PROCESS;



b2v_inst97 : lpm_ff5
PORT MAP(clock => DDRCLK(2),
		 data => SR_VDMP,
		 q => VDMP);


b2v_sr0 : lpm_shiftreg0
PORT MAP(load => SYNTHESIZED_WIRE_64,
		 clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 shiftin => SYNTHESIZED_WIRE_49,
		 data => FIFO_D(127 DOWNTO 112),
		 shiftout => CLUT_ADR(0));


b2v_sr1 : lpm_shiftreg0
PORT MAP(load => SYNTHESIZED_WIRE_64,
		 clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 shiftin => SYNTHESIZED_WIRE_50,
		 data => FIFO_D(111 DOWNTO 96),
		 shiftout => CLUT_ADR1A);


b2v_sr2 : lpm_shiftreg0
PORT MAP(load => SYNTHESIZED_WIRE_64,
		 clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 shiftin => SYNTHESIZED_WIRE_51,
		 data => FIFO_D(95 DOWNTO 80),
		 shiftout => CLUT_ADR2A);


b2v_sr3 : lpm_shiftreg0
PORT MAP(load => SYNTHESIZED_WIRE_64,
		 clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 shiftin => SYNTHESIZED_WIRE_52,
		 data => FIFO_D(79 DOWNTO 64),
		 shiftout => CLUT_ADR3A);


b2v_sr4 : lpm_shiftreg0
PORT MAP(load => SYNTHESIZED_WIRE_64,
		 clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 shiftin => SYNTHESIZED_WIRE_53,
		 data => FIFO_D(63 DOWNTO 48),
		 shiftout => CLUT_ADR4A);


b2v_sr5 : lpm_shiftreg0
PORT MAP(load => SYNTHESIZED_WIRE_64,
		 clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 shiftin => SYNTHESIZED_WIRE_54,
		 data => FIFO_D(47 DOWNTO 32),
		 shiftout => CLUT_ADR5A);


b2v_sr6 : lpm_shiftreg0
PORT MAP(load => SYNTHESIZED_WIRE_64,
		 clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 shiftin => CLUT_ADR7A,
		 data => FIFO_D(31 DOWNTO 16),
		 shiftout => CLUT_ADR6A);


b2v_sr7 : lpm_shiftreg0
PORT MAP(load => SYNTHESIZED_WIRE_64,
		 clock => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 shiftin => CLUT_ADR(0),
		 data => FIFO_D(15 DOWNTO 0),
		 shiftout => CLUT_ADR7A);


b2v_ST_CLUT_BLUE : altdpram0
PORT MAP(wren_a => ST_CLUT_WR(1),
		 wren_b => SYNTHESIZED_WIRE_55,
		 clock_a => MAIN_CLK,
		 clock_b => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 address_a => FB_ADR(4 DOWNTO 1),
		 address_b => CLUT_ADR(3 DOWNTO 0),
		 data_a => FB_AD(18 DOWNTO 16),
		 q_a => SYNTHESIZED_WIRE_34,
		 q_b => CCS(7 DOWNTO 5));


b2v_ST_CLUT_GREEN : altdpram0
PORT MAP(wren_a => ST_CLUT_WR(1),
		 wren_b => SYNTHESIZED_WIRE_56,
		 clock_a => MAIN_CLK,
		 clock_b => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 address_a => FB_ADR(4 DOWNTO 1),
		 address_b => CLUT_ADR(3 DOWNTO 0),
		 data_a => FB_AD(22 DOWNTO 20),
		 q_a => SYNTHESIZED_WIRE_31,
		 q_b => CCS(15 DOWNTO 13));


b2v_ST_CLUT_RED : altdpram0
PORT MAP(wren_a => ST_CLUT_WR(0),
		 wren_b => SYNTHESIZED_WIRE_57,
		 clock_a => MAIN_CLK,
		 clock_b => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 address_a => FB_ADR(4 DOWNTO 1),
		 address_b => CLUT_ADR(3 DOWNTO 0),
		 data_a => FB_AD(26 DOWNTO 24),
		 q_a => SYNTHESIZED_WIRE_29,
		 q_b => CCS(23 DOWNTO 21));


b2v_VIDEO_MOD_MUX_CLUTCTR : video_mod_mux_clutctr
PORT MAP(nRSTO => nRSTO,
		 MAIN_CLK => MAIN_CLK,
		 nFB_CS1 => nFB_CS1,
		 nFB_CS2 => nFB_CS2,
		 nFB_CS3 => nFB_CS3,
		 nFB_WR => nFB_WR,
		 nFB_OE => nFB_OE,
		 FB_SIZE0 => FB_SIZE0,
		 FB_SIZE1 => FB_SIZE1,
		 nFB_BURST => nFB_BURST,
		 CLK33M => CLK33M,
		 CLK25M => CLK25M,
		 BLITTER_RUN => BLITTER_RUN,
		 CLK_VIDEO => CLK_VIDEO,
		 VR_BUSY => VR_BUSY,
		 FB_AD => FB_AD,
		 FB_ADR => FB_ADR,
		 VR_D => VR_D,
		 COLOR8 => COLOR8,
		 ACP_CLUT_RD => ACP_CLUT_RD,
		 COLOR1 => COLOR1,
		 FALCON_CLUT_RDH => FALCON_CLUT_RDH,
		 FALCON_CLUT_RDL => FALCON_CLUT_RDL,
		 ST_CLUT_RD => ST_CLUT_RD,
		 HSYNC => HSYNC,
		 VSYNC => VSYNC,
		 nBLANK => nBLANK,
		 nSYNC => nSYNC,
		 nPD_VGA => nPD_VGA,
		 FIFO_RDE => FIFO_RDE,
		 COLOR2 => COLOR2,
		 COLOR4 => COLOR4,
		 PIXEL_CLK => PIXEL_CLK_ALTERA_SYNTHESIZED,
		 BLITTER_ON => BLITTER_ON,
		 VIDEO_MOD_TA => VIDEO_MOD_TA,
		 INTER_ZEI => INTER_ZEI,
		 DOP_FIFO_CLR => DOP_FIFO_CLR,
		 VIDEO_RECONFIG => VIDEO_RECONFIG,
		 VR_WR => VR_WR,
		 VR_RD => VR_RD,
		 CLR_FIFO => CLR_FIFO,
		 ACP_CLUT_WR => ACP_CLUT_WR,
		 CCR => CCR,
		 CCSEL => CCSEL,
		 CLUT_MUX_ADR => CLUT_MUX_ADR,
		 CLUT_OFF => CLUT_OFF,
		 FALCON_CLUT_WR => FALCON_CLUT_WR,
		 ST_CLUT_WR => ST_CLUT_WR,
		 VIDEO_RAM_CTR => VIDEO_RAM_CTR);

PIXEL_CLK <= PIXEL_CLK_ALTERA_SYNTHESIZED;

END bdf_type;